`timescale 1ns / 1ps
`default_nettype none
`define CODE {OPcode,Fun3,Fun12}
`define CONTROL {ALU_Control, ALUSrc_B, Branch, Jump, MemRead, MemtoReg, MemWrite, RegWrite, ill_inst, mret, ecall}

module SCPU_ctrl(input wire [6:0] OPcode,
                 input wire [2:0] Fun3,
                 input wire [11:0] Fun12,
                 output reg [3:0] ALU_Control,
                 output reg ALUSrc_B,
                 output reg [1:0] Branch,
                 output reg [1:0] Jump,
                 output reg MemRead,
                 output reg [1:0] MemtoReg,
                 output reg MemWrite,
                 output reg RegWrite,
                 output reg ill_inst,
                 output reg mret,
                 output reg ecall);
    
    
    always @(*) begin
        casez(`CODE)
            22'b0110011_000_0000000_?????: `CONTROL = 17'b00100_0000_00001_000; //add
            22'b0110011_000_0100000_?????: `CONTROL = 17'b01100_0000_00001_000; //sub
            22'b0110011_100_0000000_?????: `CONTROL = 17'b00110_0000_00001_000; //xor
            22'b0110011_110_0000000_?????: `CONTROL = 17'b00010_0000_00001_000; //or
            22'b0110011_111_0000000_?????: `CONTROL = 17'b00000_0000_00001_000; //and
            22'b0110011_001_0000000_?????: `CONTROL = 17'b01000_0000_00001_000; //sll
            22'b0110011_101_0000000_?????: `CONTROL = 17'b01010_0000_00001_000; //srl
            22'b0110011_101_0100000_?????: `CONTROL = 17'b10000_0000_00001_000; //sra
            22'b0110011_010_0000000_?????: `CONTROL = 17'b01110_0000_00001_000; //slt
            22'b0110011_011_0000000_?????: `CONTROL = 17'b10010_0000_00001_000; //sltu
            22'b0010011_000_???????_?????: `CONTROL = 17'b00101_0000_00001_000; //addi
            22'b0010011_100_???????_?????: `CONTROL = 17'b00111_0000_00001_000; //xori
            22'b0010011_110_???????_?????: `CONTROL = 17'b00011_0000_00001_000; //ori
            22'b0010011_111_???????_?????: `CONTROL = 17'b00001_0000_00001_000; //andi
            22'b0010011_001_0000000_?????: `CONTROL = 17'b01001_0000_00001_000; //slli
            22'b0010011_101_0000000_?????: `CONTROL = 17'b01011_0000_00001_000; //srli
            22'b0010011_101_0100000_?????: `CONTROL = 17'b10001_0000_00001_000; //srai
            22'b0010011_010_???????_?????: `CONTROL = 17'b01111_0000_00001_000; //slti
            22'b0010011_011_???????_?????: `CONTROL = 17'b10011_0000_00001_000; //sltiu
            22'b0000011_000_???????_?????: `CONTROL = 17'b00101_0000_10101_000; //lb
            22'b0000011_001_???????_?????: `CONTROL = 17'b00101_0000_10101_000; //lh
            22'b0000011_010_???????_?????: `CONTROL = 17'b00101_0000_10101_000; //lw
            22'b0000011_100_???????_?????: `CONTROL = 17'b00101_0000_10101_000; //lbu
            22'b0000011_101_???????_?????: `CONTROL = 17'b00101_0000_10101_000; //lhu
            22'b0100011_000_???????_?????: `CONTROL = 17'b00101_0000_00010_000; //sb
            22'b0100011_001_???????_?????: `CONTROL = 17'b00101_0000_00010_000; //sh
            22'b0100011_010_???????_?????: `CONTROL = 17'b00101_0000_00010_000; //sw
            22'b1100011_000_???????_?????: `CONTROL = 17'b01100_1100_00000_000; //beq
            22'b1100011_001_???????_?????: `CONTROL = 17'b01100_1000_00000_000; //bne
            22'b1100011_100_???????_?????: `CONTROL = 17'b01110_1000_00000_000; //blt
            22'b1100011_101_???????_?????: `CONTROL = 17'b01110_1100_00000_000; //bge
            22'b1100011_110_???????_?????: `CONTROL = 17'b10010_1000_00000_000; //bltu
            22'b1100011_111_???????_?????: `CONTROL = 17'b10010_1100_00000_000; //bgeu
            22'b1101111_???_???????_?????: `CONTROL = 17'b11110_0001_01001_000; //jal
            22'b1100111_000_???????_?????: `CONTROL = 17'b11110_0010_01001_000; //jalr
            22'b0110111_???_???????_?????: `CONTROL = 17'b11110_0000_11101_000; //lui
            22'b0010111_???_???????_?????: `CONTROL = 17'b11110_0000_01101_000; //auipc
            22'b1110011_000_0000000_00000: `CONTROL = 17'b11110_0000_00000_001; //ecall
            22'b1110011_000_0000000_00001: `CONTROL = 17'b11110_0000_00000_001; //ebreak
            22'b1110011_000_0011000_00010: `CONTROL = 17'b11110_0000_00000_010; //mret
            default: `CONTROL                       = 17'b11110_0000_00000_100; //ILLEGAL
        endcase
    end
    
endmodule
